*** SPICE deck for cell control_logic_test{sch} from library ese370project2
*** Created on Sat Dec 02, 2017 13:02:05
*** Last revised on Sun Dec 03, 2017 00:34:49
*** Written on Sun Dec 03, 2017 00:35:56 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 22nm_HP.pm

*** SUBCIRCUIT ese370project2__buffer FROM CELL buffer{sch}
.SUBCKT ese370project2__buffer ground in o power
Mnmos@0 net@13 in ground ground N L=0.022U W=0.022U
Mnmos@1 o net@13 ground ground N L=0.022U W=0.022U
Mpmos@0 power in net@13 power P L=0.022U W=0.022U
Mpmos@1 power net@13 o power P L=0.022U W=0.022U
.ENDS ese370project2__buffer

*** SUBCIRCUIT ese370project2__inv FROM CELL inv{sch}
.SUBCKT ese370project2__inv ground in o power
Mnmos@0 o in ground ground N L=0.022U W=0.022U
Mpmos@0 power in o power P L=0.022U W=0.022U
.ENDS ese370project2__inv

*** SUBCIRCUIT ese370project2__nor2_clock FROM CELL nor2_clock{sch}
.SUBCKT ese370project2__nor2_clock A B Ground Out Power
Mnmos@0 Out A Ground Ground N L=0.022U W=0.352U
Mnmos@1 Out B Ground Ground N L=0.022U W=0.352U
Mpmos@0 Power A net@0 Power P L=0.022U W=0.352U
Mpmos@1 net@0 B Out Power P L=0.022U W=0.352U
.ENDS ese370project2__nor2_clock

*** SUBCIRCUIT ese370project2__clock_gen FROM CELL clock_gen{sch}
.SUBCKT ese370project2__clock_gen clk clk_n ground in power
Mnmos@0 net@90 net@38 ground ground N L=0.022U W=0.704U
Mnmos@1 clk net@90 ground ground N L=0.022U W=1.408U
Mnmos@2 net@113 net@41 ground ground N L=0.022U W=0.704U
Mnmos@3 clk_n net@113 ground ground N L=0.022U W=1.408U
Mpmos@0 power net@38 net@90 power P L=0.022U W=0.704U
Mpmos@1 power net@90 clk power P L=0.022U W=1.408U
Mpmos@2 power net@41 net@113 power P L=0.022U W=0.704U
Mpmos@3 power net@113 clk_n power P L=0.022U W=1.408U
Xbuffer@0 ground in net@74 power ese370project2__buffer
Xinv@0 ground in net@67 power ese370project2__inv
Xnor2_clo@0 net@67 net@41 ground net@38 power ese370project2__nor2_clock
Xnor2_clo@1 net@38 net@74 ground net@41 power ese370project2__nor2_clock
.ENDS ese370project2__clock_gen

*** SUBCIRCUIT ese370project2__nand2 FROM CELL nand2{sch}
.SUBCKT ese370project2__nand2 A B Ground O Power
Mnmos@0 O A net@36 Ground N L=0.022U W=0.022U
Mnmos@1 net@36 B Ground Ground N L=0.022U W=0.022U
Mpmos@0 Power A O Power P L=0.022U W=0.022U
Mpmos@1 Power B O Power P L=0.022U W=0.022U
.ENDS ese370project2__nand2

*** SUBCIRCUIT ese370project2__gate_based_latch FROM CELL gate_based_latch{sch}
.SUBCKT ese370project2__gate_based_latch Ground In Out Phi Power
Xinv@1 Ground Phi net@22 Power ese370project2__inv
Xnand2@0 In Phi Ground net@10 Power ese370project2__nand2
Xnand2@1 net@22 Out Ground net@6 Power ese370project2__nand2
Xnand2@2 net@10 net@6 Ground Out Power ese370project2__nand2
.ENDS ese370project2__gate_based_latch

*** SUBCIRCUIT ese370project2__gate_based_register FROM CELL gate_based_register{sch}
.SUBCKT ese370project2__gate_based_register Clk0 Clk1 Ground In Out Out_n Power
Xgate_bas@0 Ground In net@0 Clk0 Power ese370project2__gate_based_latch
Xgate_bas@1 Ground net@0 Out Clk1 Power ese370project2__gate_based_latch
Xinv@0 Ground Out Out_n Power ese370project2__inv
.ENDS ese370project2__gate_based_register

*** SUBCIRCUIT ese370project2__clock_box FROM CELL clock_box{sch}
.SUBCKT ese370project2__clock_box _1Ghz _1Ghz_n _500Mhz _500Mhz_n gnd in pwr
Xclock_ge@0 _500Mhz _500Mhz_n gnd net@11 pwr ese370project2__clock_gen
Xclock_ge@1 _1Ghz _1Ghz_n gnd in pwr ese370project2__clock_gen
Xgate_bas@0 net@43 in gnd net@0 net@11 net@0 pwr ese370project2__gate_based_register
Xinv@0 gnd in net@43 pwr ese370project2__inv
.ENDS ese370project2__clock_box

*** SUBCIRCUIT ese370project2__nor4 FROM CELL nor4{sch}
.SUBCKT ese370project2__nor4 A B C D Ground Out Power
Mnmos@0 Out A Ground Ground N L=0.022U W=0.022U
Mnmos@1 Out B Ground Ground N L=0.022U W=0.022U
Mnmos@2 Out C Ground Ground N L=0.022U W=0.022U
Mnmos@3 Out D Ground Ground N L=0.022U W=0.022U
Mpmos@0 net@28 C net@0 Power P L=0.022U W=0.022U
Mpmos@1 net@0 D Out Power P L=0.022U W=0.022U
Mpmos@2 Power A net@27 Power P L=0.022U W=0.022U
Mpmos@3 net@27 B net@28 Power P L=0.022U W=0.022U
.ENDS ese370project2__nor4

*** SUBCIRCUIT ese370project2__xor2 FROM CELL xor2{sch}
.SUBCKT ese370project2__xor2 A B gnd out pwr
Xnand2@0 A B gnd net@21 pwr ese370project2__nand2
Xnand2@1 net@21 B gnd net@0 pwr ese370project2__nand2
Xnand2@2 A net@21 gnd net@3 pwr ese370project2__nand2
Xnand2@3 net@3 net@0 gnd out pwr ese370project2__nand2
.ENDS ese370project2__xor2

*** SUBCIRCUIT ese370project2__comparator FROM CELL comparator{sch}
.SUBCKT ese370project2__comparator a0 a1 a2 a3 b0 b1 b2 b3 gnd out pwr
Xnor4@0 net@51 net@48 net@45 net@42 gnd out pwr ese370project2__nor4
Xxor2@0 a0 b0 gnd net@51 pwr ese370project2__xor2
Xxor2@1 a1 b1 gnd net@48 pwr ese370project2__xor2
Xxor2@2 a2 b2 gnd net@45 pwr ese370project2__xor2
Xxor2@3 a3 b3 gnd net@42 pwr ese370project2__xor2
.ENDS ese370project2__comparator

*** SUBCIRCUIT ese370project2__counter FROM CELL counter{sch}
.SUBCKT ese370project2__counter c0 c1 c2 c3 clk clk_n gnd pwr
Xgate_bas@0 clk clk_n gnd net@0 c0 net@0 pwr ese370project2__gate_based_register
Xgate_bas@1 c0 net@0 gnd net@51 c1 net@51 pwr ese370project2__gate_based_register
Xgate_bas@3 c1 net@51 gnd net@81 c2 net@81 pwr ese370project2__gate_based_register
Xgate_bas@5 c2 net@81 gnd net@99 c3 net@99 pwr ese370project2__gate_based_register
.ENDS ese370project2__counter

*** SUBCIRCUIT ese370project2__nand3 FROM CELL nand3{sch}
.SUBCKT ese370project2__nand3 A B C gnd out pwr
Mnmos@0 out A net@9 gnd N L=0.022U W=0.022U
Mnmos@1 net@9 B net@10 gnd N L=0.022U W=0.022U
Mnmos@2 net@10 C gnd gnd N L=0.022U W=0.022U
Mpmos@0 pwr C out pwr P L=0.022U W=0.022U
Mpmos@1 pwr B out pwr P L=0.022U W=0.022U
Mpmos@2 pwr A out pwr P L=0.022U W=0.022U
.ENDS ese370project2__nand3

*** SUBCIRCUIT ese370project2__bitslice FROM CELL bitslice{sch}
.SUBCKT ese370project2__bitslice A B Cin Cout gnd pwr S
Xnand2@0 A Cin gnd net@5 pwr ese370project2__nand2
Xnand2@1 A B gnd net@107 pwr ese370project2__nand2
Xnand2@2 B Cin gnd net@1 pwr ese370project2__nand2
Xnand3@0 net@5 net@107 net@1 gnd Cout pwr ese370project2__nand3
Xxor2@0 B A gnd net@9 pwr ese370project2__xor2
Xxor2@1 net@9 Cin gnd S pwr ese370project2__xor2
.ENDS ese370project2__bitslice

*** SUBCIRCUIT ese370project2__four_adder FROM CELL four_adder{sch}
.SUBCKT ese370project2__four_adder a0 a1 a2 a3 b0 b1 b2 b3 gnd pwr s0 s1 s2 s3
Xbitslice@0 a1 b1 net@20 net@26 gnd pwr s1 ese370project2__bitslice
Xbitslice@1 a2 b2 net@26 net@31 gnd pwr s2 ese370project2__bitslice
Xbitslice@2 a3 b3 net@31 net@41 gnd pwr s3 ese370project2__bitslice
Xbitslice@3 a0 b0 gnd net@20 gnd pwr s0 ese370project2__bitslice
.ENDS ese370project2__four_adder

*** SUBCIRCUIT ese370project2__counter_logic FROM CELL counter_logic{sch}
.SUBCKT ese370project2__counter_logic empty full ground head head0 head1 head2 head3 power tail tail0 tail1 tail2 tail3
Xcomparat@0 net@226 net@225 net@182 net@184 tail0 tail1 tail2 tail3 ground full power ese370project2__comparator
Xcomparat@1 head0 head1 head2 head3 tail0 tail1 tail2 tail3 ground empty power ese370project2__comparator
Xcounter@0 head0 head1 head2 head3 head net@52 ground power ese370project2__counter
Xcounter@1 tail0 tail1 tail2 tail3 tail net@58 ground power ese370project2__counter
Xfour_add@0 head0 head1 head2 head3 power ground ground ground ground power net@226 net@225 net@182 net@184 ese370project2__four_adder
Xinv@0 ground head net@52 power ese370project2__inv
Xinv@1 ground tail net@58 power ese370project2__inv
.ENDS ese370project2__counter_logic

*** SUBCIRCUIT ese370project2__nor2 FROM CELL nor2{sch}
.SUBCKT ese370project2__nor2 A B Ground Out Power
Mnmos@0 Out A Ground Ground N L=0.022U W=0.022U
Mnmos@1 Out B Ground Ground N L=0.022U W=0.022U
Mpmos@0 Power A net@0 Power P L=0.022U W=0.022U
Mpmos@1 net@0 B Out Power P L=0.022U W=0.022U
.ENDS ese370project2__nor2

*** SUBCIRCUIT ese370project2__control_logic FROM CELL control_logic{sch}
.SUBCKT ese370project2__control_logic deq empty enq full ghz gnd head0 head1 head2 head3 mhz pwr read tail0 tail1 tail2 tail3 write
Mnmos@0 net@287 net@130 gnd gnd N L=0.022U W=0.088U
Mnmos@1 read net@287 gnd gnd N L=0.022U W=0.352U
Mnmos@2 net@310 net@127 gnd gnd N L=0.022U W=0.088U
Mnmos@3 write net@310 gnd gnd N L=0.022U W=0.352U
Mpmos@0 pwr net@130 net@287 pwr P L=0.022U W=0.088U
Mpmos@1 pwr net@287 read pwr P L=0.022U W=0.352U
Mpmos@2 pwr net@127 net@310 pwr P L=0.022U W=0.088U
Mpmos@3 pwr net@310 write pwr P L=0.022U W=0.352U
Xcounter_@0 empty full gnd net@127 head0 head1 head2 head3 pwr net@130 tail0 tail1 tail2 tail3 ese370project2__counter_logic
Xinv@0 gnd net@188 net@130 pwr ese370project2__inv
Xinv@1 gnd net@230 net@127 pwr ese370project2__inv
Xinv@3 gnd net@34 net@38 pwr ese370project2__inv
Xinv@4 gnd ghz net@91 pwr ese370project2__inv
Xinv@8 gnd empty net@200 pwr ese370project2__inv
Xinv@9 gnd full net@175 pwr ese370project2__inv
Xnand2@3 net@91 mhz gnd net@34 pwr ese370project2__nand2
Xnand3@2 enq net@175 net@38 gnd net@230 pwr ese370project2__nand3
Xnand3@3 net@82 net@200 deq gnd net@188 pwr ese370project2__nand3
Xnor2@1 ghz mhz gnd net@82 pwr ese370project2__nor2
.ENDS ese370project2__control_logic

.global gnd vdd

*** TOP LEVEL CELL: control_logic_test{sch}
VVPWL@0 deq gnd pwl (0ns 0 1.6ns 0 1.61ns 0.8 2ns 0.8 2.01ns 0) DC 0V AC 0V 0
VVPWL@1 enq gnd pwl (0ns 0.8 0.99ns 0.8 1ns 0 2ns 0 2.01 0.8) DC 0V AC 0V 0
VVPulse@0 net@29 gnd pulse (0 0.8V 0ns 10ps 10ps 0.5ns 1ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xclock_bo@0 ghz clock_bo@0_1Ghz_n mhz clock_bo@0_500Mhz_n gnd net@29 vdd ese370project2__clock_box
Xcontrol_@0 deq empty enq full ghz gnd head0 head1 head2 head3 mhz vdd read tail0 tail1 tail2 tail3 write ese370project2__control_logic
.END
