*** SPICE deck for cell tristate_buffer_test{sch} from library ese370project2
*** Created on Sun Nov 19, 2017 18:09:32
*** Last revised on Sun Nov 19, 2017 18:12:46
*** Written on Sun Nov 19, 2017 18:12:55 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 22nm_HP.pm

*** SUBCIRCUIT ese370project2__tristate_buffer FROM CELL tristate_buffer{sch}
.SUBCKT ese370project2__tristate_buffer en ground in out power
Mnmos@0 net@1 net@4 ground ground N L=0.022U W=0.022U
Mnmos@1 out en net@1 ground N L=0.022U W=0.022U
Mnmos@2 net@4 in ground ground N L=0.022U W=0.022U
Mpmos@0 power net@4 net@1 power P L=0.022U W=0.022U
Mpmos@1 power in net@4 power P L=0.022U W=0.022U
.ENDS ese370project2__tristate_buffer

.global gnd vdd

*** TOP LEVEL CELL: tristate_buffer_test{sch}
VVPulse@0 net_en gnd pulse (0 0.8V 0ns 10ps 10ps 1ns 2ns) DC 0V AC 0V 0
VVPulse@1 net_in gnd pulse (0 0.8V 0ns 10ps 10ps 500ps 1ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xtristate@0 net_en gnd net_in net_out vdd ese370project2__tristate_buffer
.END
