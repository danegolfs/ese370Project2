*** SPICE deck for cell sense_amp_test{sch} from library ese370project2
*** Created on Sun Nov 19, 2017 18:09:18
*** Last revised on Sun Nov 19, 2017 19:24:55
*** Written on Sun Nov 19, 2017 19:25:01 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 22nm_HP.pm

*** SUBCIRCUIT ese370project2__sense_amp FROM CELL sense_amp{sch}
.SUBCKT ese370project2__sense_amp en ground in n_in out power
Mnmos@1 net@20 n_in out ground N L=0.022U W=0.022U
Mnmos@2 net@20 en ground ground N L=0.022U W=0.022U
Mnmos@3 net@8 in net@20 ground N L=0.022U W=0.022U
Mpmos@0 net@8 net@8 power power P L=0.022U W=0.022U
Mpmos@1 power net@8 out power P L=0.022U W=0.022U
.ENDS ese370project2__sense_amp

.global gnd vdd

*** TOP LEVEL CELL: sense_amp_test{sch}
VVPWL@0 net_in gnd pwl (0ns 0 500ps 0.8 1ns 0 1500ps 0.8 2ns 0) DC 0V AC 0V 0
VVPulse@0 net_en gnd pulse (0 0.8V 0ns 10ps 10ps 1ns 2ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
VV_Generi@1 net_n_in gnd DC 0.4 AC 0
Xsense_am@0 net_en gnd net_in net_n_in net_out vdd ese370project2__sense_amp
.END
