*** SPICE deck for cell clock_box_test{sch} from library ese370project2
*** Created on Mon Dec 04, 2017 18:33:01
*** Last revised on Mon Dec 04, 2017 18:35:20
*** Written on Mon Dec 04, 2017 18:35:24 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 22nm_HP.pm

*** SUBCIRCUIT ese370project2__buffer FROM CELL buffer{sch}
.SUBCKT ese370project2__buffer ground in o power
Mnmos@0 net@13 in ground ground N L=0.022U W=0.022U
Mnmos@1 o net@13 ground ground N L=0.022U W=0.022U
Mpmos@0 power in net@13 power P L=0.022U W=0.022U
Mpmos@1 power net@13 o power P L=0.022U W=0.022U
.ENDS ese370project2__buffer

*** SUBCIRCUIT ese370project2__inv FROM CELL inv{sch}
.SUBCKT ese370project2__inv ground in o power
Mnmos@0 o in ground ground N L=0.022U W=0.022U
Mpmos@0 power in o power P L=0.022U W=0.022U
.ENDS ese370project2__inv

*** SUBCIRCUIT ese370project2__nor2_clock FROM CELL nor2_clock{sch}
.SUBCKT ese370project2__nor2_clock A B Ground Out Power
Mnmos@0 Out A Ground Ground N L=0.022U W=0.352U
Mnmos@1 Out B Ground Ground N L=0.022U W=0.352U
Mpmos@0 Power A net@0 Power P L=0.022U W=0.352U
Mpmos@1 net@0 B Out Power P L=0.022U W=0.352U
.ENDS ese370project2__nor2_clock

*** SUBCIRCUIT ese370project2__clock_gen FROM CELL clock_gen{sch}
.SUBCKT ese370project2__clock_gen clk clk_n ground in power
Mnmos@0 net@90 net@38 ground ground N L=0.022U W=0.704U
Mnmos@1 clk net@90 ground ground N L=0.022U W=1.408U
Mnmos@2 net@113 net@41 ground ground N L=0.022U W=0.704U
Mnmos@3 clk_n net@113 ground ground N L=0.022U W=1.408U
Mpmos@0 power net@38 net@90 power P L=0.022U W=0.704U
Mpmos@1 power net@90 clk power P L=0.022U W=1.408U
Mpmos@2 power net@41 net@113 power P L=0.022U W=0.704U
Mpmos@3 power net@113 clk_n power P L=0.022U W=1.408U
Xbuffer@0 ground in net@74 power ese370project2__buffer
Xinv@0 ground in net@67 power ese370project2__inv
Xnor2_clo@0 net@67 net@41 ground net@38 power ese370project2__nor2_clock
Xnor2_clo@1 net@38 net@74 ground net@41 power ese370project2__nor2_clock
.ENDS ese370project2__clock_gen

*** SUBCIRCUIT ese370project2__nand2 FROM CELL nand2{sch}
.SUBCKT ese370project2__nand2 A B Ground O Power
Mnmos@0 O A net@36 Ground N L=0.022U W=0.022U
Mnmos@1 net@36 B Ground Ground N L=0.022U W=0.022U
Mpmos@0 Power A O Power P L=0.022U W=0.022U
Mpmos@1 Power B O Power P L=0.022U W=0.022U
.ENDS ese370project2__nand2

*** SUBCIRCUIT ese370project2__gate_based_latch FROM CELL gate_based_latch{sch}
.SUBCKT ese370project2__gate_based_latch Ground In Out Phi Power
Xinv@1 Ground Phi net@22 Power ese370project2__inv
Xnand2@0 In Phi Ground net@10 Power ese370project2__nand2
Xnand2@1 net@22 Out Ground net@6 Power ese370project2__nand2
Xnand2@2 net@10 net@6 Ground Out Power ese370project2__nand2
.ENDS ese370project2__gate_based_latch

*** SUBCIRCUIT ese370project2__gate_based_register FROM CELL gate_based_register{sch}
.SUBCKT ese370project2__gate_based_register Clk0 Clk1 Ground In Out Out_n Power
Xgate_bas@0 Ground In net@0 Clk0 Power ese370project2__gate_based_latch
Xgate_bas@1 Ground net@0 Out Clk1 Power ese370project2__gate_based_latch
Xinv@0 Ground Out Out_n Power ese370project2__inv
.ENDS ese370project2__gate_based_register

*** SUBCIRCUIT ese370project2__clock_box FROM CELL clock_box{sch}
.SUBCKT ese370project2__clock_box _1Ghz _1Ghz_n _500Mhz _500Mhz_n gnd in pwr
Xclock_ge@0 _500Mhz _500Mhz_n gnd net@11 pwr ese370project2__clock_gen
Xclock_ge@1 _1Ghz _1Ghz_n gnd in pwr ese370project2__clock_gen
Xgate_bas@0 net@43 in gnd net@0 net@11 net@0 pwr ese370project2__gate_based_register
Xinv@0 gnd in net@43 pwr ese370project2__inv
.ENDS ese370project2__clock_box

.global gnd vdd

*** TOP LEVEL CELL: clock_box_test{sch}
VVPulse@0 net@2 gnd pulse (0 0.8V 0ns 10ps 10ps 0.5ns 1ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xclock_bo@0 ghz ghz_n mhz mhz_n gnd net@2 vdd ese370project2__clock_box
.END
