*** SPICE deck for cell test_transistor_capacitance{sch} from library ese370project2
*** Created on Tue Nov 21, 2017 13:56:59
*** Last revised on Tue Nov 21, 2017 14:05:55
*** Written on Tue Nov 21, 2017 14:06:00 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 22nm_HP.pm

.global gnd vdd

*** TOP LEVEL CELL: test_transistor_capacitance{sch}
Mnmos@0 gnd net_out1 gnd gnd N L=0.022U W=0.022U
Mnmos@1 net_out1 gnd gnd gnd N L=0.022U W=0.022U
Mnmos@2 gnd net_out2 gnd gnd N L=0.022U W=0.044U
Mnmos@4 net_out3 gnd gnd gnd N L=0.022U W=0.044U
Mnmos@6 net_out1 net_in gnd gnd N L=0.022U W=0.022U
Mnmos@7 net_out2 net_in gnd gnd N L=0.022U W=0.022U
Mnmos@8 net_out3 net_in gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd net_in net_out1 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net_in net_out2 vdd P L=0.022U W=0.022U
Mpmos@2 vdd net_in net_out3 vdd P L=0.022U W=0.022U
VVPulse@0 net_in gnd pulse (0 0.8V 0ns 1fs 1fs 1ns 2ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
.END
