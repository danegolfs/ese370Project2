*** SPICE deck for cell tristate_buffer_test{sch} from library ese370project2
*** Created on Sun Nov 19, 2017 18:09:32
*** Last revised on Mon Dec 04, 2017 18:55:56
*** Written on Mon Dec 04, 2017 18:56:19 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 22nm_HP.pm

*** SUBCIRCUIT ese370project2__tristate_buffer_min_size FROM CELL tristate_buffer_min_size{sch}
.SUBCKT ese370project2__tristate_buffer_min_size en ground in out power
Mnmos@0 out net@11 net@31 ground N L=0.022U W=0.022U
Mnmos@1 net@11 in ground ground N L=0.022U W=0.022U
Mnmos@2 net@31 en ground ground N L=0.022U W=0.022U
Mnmos@3 net@1 en ground ground N L=0.022U W=0.022U
Mpmos@0 net@29 net@11 out power P L=0.022U W=0.022U
Mpmos@1 power in net@11 power P L=0.022U W=0.022U
Mpmos@2 power net@1 net@29 power P L=0.022U W=0.022U
Mpmos@3 power en net@1 power P L=0.022U W=0.022U
.ENDS ese370project2__tristate_buffer_min_size

.global gnd vdd

*** TOP LEVEL CELL: tristate_buffer_test{sch}
Mnmos@0 net@13 net_out net@13 gnd N L=0.022U W=0.088U
VVPulse@0 net_en gnd pulse (0 0.8V 0ns 10ps 10ps 1ns 2ns) DC 0V AC 0V 0
VVPulse@1 net_in gnd pulse (0 0.8V 0ns 10ps 10ps 500ps 1ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xtristate@1 net_en gnd net_in net_out vdd ese370project2__tristate_buffer_min_size
.END
