*** SPICE deck for cell celltest{sch} from library ese370project2
*** Created on Sat Nov 18, 2017 14:46:32
*** Last revised on Sun Nov 19, 2017 13:03:30
*** Written on Sun Nov 19, 2017 13:04:20 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 22nm_HP.pm

*** SUBCIRCUIT ese370project2__5TCell FROM CELL 5TCell{sch}
.SUBCKT ese370project2__5TCell A bitline enable ground power
Mnmos@2 bitline enable A ground N L=0.022U W=0.022U
Mnmos@3 net@10 A ground ground N L=0.022U W=0.022U
Mnmos@4 A net@10 ground ground N L=0.022U W=0.022U
Mpmos@2 power A net@10 power P L=0.022U W=0.022U
Mpmos@3 power net@10 A power P L=0.022U W=0.022U
.ENDS ese370project2__5TCell

.global gnd vdd

*** TOP LEVEL CELL: celltest{sch}
Mnmos@0 net_BL net_drive_enable net_drive gnd N L=0.022U W=0.022U
X_5TCell@0 net_A net_BL net_WL gnd vdd ese370project2__5TCell
VV_Generi@0 vdd gnd DC 0.8 AC 0
Vdrive net_drive gnd pwl (0ns 0 1.99ns 0 2.0ns 0.8V 3.99ns 0.8V 4.0ns 0 4.99ns 0 5.0ns 0.4V 5.49ns 0.4V 5.50ns 0 7.98ns 0 ) DC 0V AC 0V 0
VdriveE net_drive_enable gnd pwl (0ns 0 1.98ns 0 1.99ns 0.8V 3.98ns 0.8V 3.99ns 0 4.98ns 0 4.99ns 0.8V 5.48ns 0.8V 5.49ns 0 7.98ns) DC 0V AC 0V 0
Venable net_WL gnd pwl (0ns 0 1.98ns 0 1.99ns 0.8V 3.98ns 0.8V 3.99ns 0 5.98ns 0 5.99ns 0.8V 7.98ns 0.8V 7.99ns 0) DC 0V AC 0V 0
.END
