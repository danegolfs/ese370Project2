*** SPICE deck for cell counter_logic_test{sch} from library ese370project2
*** Created on Sat Dec 02, 2017 13:01:14
*** Last revised on Sun Dec 03, 2017 14:16:00
*** Written on Mon Dec 04, 2017 19:36:31 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 22nm_HP.pm

*** SUBCIRCUIT ese370project2__nor4 FROM CELL nor4{sch}
.SUBCKT ese370project2__nor4 A B C D Ground Out Power
Mnmos@0 Out A Ground Ground N L=0.022U W=0.022U
Mnmos@1 Out B Ground Ground N L=0.022U W=0.022U
Mnmos@2 Out C Ground Ground N L=0.022U W=0.022U
Mnmos@3 Out D Ground Ground N L=0.022U W=0.022U
Mpmos@0 net@28 C net@0 Power P L=0.022U W=0.022U
Mpmos@1 net@0 D Out Power P L=0.022U W=0.022U
Mpmos@2 Power A net@27 Power P L=0.022U W=0.022U
Mpmos@3 net@27 B net@28 Power P L=0.022U W=0.022U
.ENDS ese370project2__nor4

*** SUBCIRCUIT ese370project2__nand2 FROM CELL nand2{sch}
.SUBCKT ese370project2__nand2 A B Ground O Power
Mnmos@0 O A net@36 Ground N L=0.022U W=0.022U
Mnmos@1 net@36 B Ground Ground N L=0.022U W=0.022U
Mpmos@0 Power A O Power P L=0.022U W=0.022U
Mpmos@1 Power B O Power P L=0.022U W=0.022U
.ENDS ese370project2__nand2

*** SUBCIRCUIT ese370project2__xor2 FROM CELL xor2{sch}
.SUBCKT ese370project2__xor2 A B gnd out pwr
Xnand2@0 A B gnd net@21 pwr ese370project2__nand2
Xnand2@1 net@21 B gnd net@0 pwr ese370project2__nand2
Xnand2@2 A net@21 gnd net@3 pwr ese370project2__nand2
Xnand2@3 net@3 net@0 gnd out pwr ese370project2__nand2
.ENDS ese370project2__xor2

*** SUBCIRCUIT ese370project2__comparator FROM CELL comparator{sch}
.SUBCKT ese370project2__comparator a0 a1 a2 a3 b0 b1 b2 b3 gnd out pwr
Xnor4@0 net@51 net@48 net@45 net@42 gnd out pwr ese370project2__nor4
Xxor2@0 a0 b0 gnd net@51 pwr ese370project2__xor2
Xxor2@1 a1 b1 gnd net@48 pwr ese370project2__xor2
Xxor2@2 a2 b2 gnd net@45 pwr ese370project2__xor2
Xxor2@3 a3 b3 gnd net@42 pwr ese370project2__xor2
.ENDS ese370project2__comparator

*** SUBCIRCUIT ese370project2__nand3 FROM CELL nand3{sch}
.SUBCKT ese370project2__nand3 A B C gnd out pwr
Mnmos@0 out A net@9 gnd N L=0.022U W=0.022U
Mnmos@1 net@9 B net@10 gnd N L=0.022U W=0.022U
Mnmos@2 net@10 C gnd gnd N L=0.022U W=0.022U
Mpmos@0 pwr C out pwr P L=0.022U W=0.022U
Mpmos@1 pwr B out pwr P L=0.022U W=0.022U
Mpmos@2 pwr A out pwr P L=0.022U W=0.022U
.ENDS ese370project2__nand3

*** SUBCIRCUIT ese370project2__bitslice FROM CELL bitslice{sch}
.SUBCKT ese370project2__bitslice A B Cin Cout gnd pwr S
Xnand2@0 A Cin gnd net@5 pwr ese370project2__nand2
Xnand2@1 A B gnd net@107 pwr ese370project2__nand2
Xnand2@2 B Cin gnd net@1 pwr ese370project2__nand2
Xnand3@0 net@5 net@107 net@1 gnd Cout pwr ese370project2__nand3
Xxor2@0 B A gnd net@9 pwr ese370project2__xor2
Xxor2@1 net@9 Cin gnd S pwr ese370project2__xor2
.ENDS ese370project2__bitslice

*** SUBCIRCUIT ese370project2__four_adder FROM CELL four_adder{sch}
.SUBCKT ese370project2__four_adder a0 a1 a2 a3 b0 b1 b2 b3 gnd pwr s0 s1 s2 s3
Xbitslice@0 a1 b1 net@20 net@26 gnd pwr s1 ese370project2__bitslice
Xbitslice@1 a2 b2 net@26 net@31 gnd pwr s2 ese370project2__bitslice
Xbitslice@2 a3 b3 net@31 net@41 gnd pwr s3 ese370project2__bitslice
Xbitslice@3 a0 b0 gnd net@20 gnd pwr s0 ese370project2__bitslice
.ENDS ese370project2__four_adder

*** SUBCIRCUIT ese370project2__inv FROM CELL inv{sch}
.SUBCKT ese370project2__inv ground in o power
Mnmos@0 o in ground ground N L=0.022U W=0.022U
Mpmos@0 power in o power P L=0.022U W=0.022U
.ENDS ese370project2__inv

*** SUBCIRCUIT ese370project2__gate_based_latch FROM CELL gate_based_latch{sch}
.SUBCKT ese370project2__gate_based_latch Ground In Out Phi Power
Xinv@1 Ground Phi net@22 Power ese370project2__inv
Xnand2@0 In Phi Ground net@10 Power ese370project2__nand2
Xnand2@1 net@22 Out Ground net@6 Power ese370project2__nand2
Xnand2@2 net@10 net@6 Ground Out Power ese370project2__nand2
.ENDS ese370project2__gate_based_latch

*** SUBCIRCUIT ese370project2__gate_based_register FROM CELL gate_based_register{sch}
.SUBCKT ese370project2__gate_based_register Clk0 Clk1 Ground In Out Out_n Power
Xgate_bas@0 Ground In net@0 Clk0 Power ese370project2__gate_based_latch
Xgate_bas@1 Ground net@0 Out Clk1 Power ese370project2__gate_based_latch
Xinv@0 Ground Out Out_n Power ese370project2__inv
.ENDS ese370project2__gate_based_register

*** SUBCIRCUIT ese370project2__register_4b FROM CELL register_4b{sch}
.SUBCKT ese370project2__register_4b clk clk_n ground in0 in1 in2 in3 out0 out1 out2 out3 power
Xgate_bas@0 clk clk_n ground in0 out0 gate_bas@0_Out_n power ese370project2__gate_based_register
Xgate_bas@1 clk clk_n ground in1 out1 gate_bas@1_Out_n power ese370project2__gate_based_register
Xgate_bas@2 clk clk_n ground in2 out2 gate_bas@2_Out_n power ese370project2__gate_based_register
Xgate_bas@3 clk clk_n ground in3 out3 gate_bas@3_Out_n power ese370project2__gate_based_register
.ENDS ese370project2__register_4b

*** SUBCIRCUIT ese370project2__counter_logic FROM CELL counter_logic{sch}
.SUBCKT ese370project2__counter_logic ground head head0 head1 head2 head3 one power sixteen tail tail0 tail1 tail2 tail3 zero
Xcomparat@0 head0 head1 head2 head3 tail0 tail1 tail2 tail3 ground zero power ese370project2__comparator
Xcomparat@1 head0 head1 head2 head3 next_tail0 next_tail1 next_tail2 next_tail3 ground one power ese370project2__comparator
Xcomparat@2 next_head0 next_head1 next_head2 next_head3 tail0 tail1 tail2 tail3 ground sixteen power ese370project2__comparator
Xfour_add@1 power ground ground ground head0 head1 head2 head3 ground power next_head0 next_head1 next_head2 next_head3 ese370project2__four_adder
Xfour_add@2 power ground ground ground tail0 tail1 tail2 tail3 ground power next_tail0 next_tail1 next_tail2 next_tail3 ese370project2__four_adder
Xinv@0 ground head net@270 power ese370project2__inv
Xinv@1 ground tail net@261 power ese370project2__inv
Xregister@0 head net@270 ground next_head0 next_head1 next_head2 next_head3 head0 head1 head2 head3 power ese370project2__register_4b
Xregister@1 tail net@261 ground next_tail0 next_tail1 next_tail2 next_tail3 tail0 tail1 tail2 tail3 power ese370project2__register_4b
.ENDS ese370project2__counter_logic

.global gnd vdd

*** TOP LEVEL CELL: counter_logic_test{sch}
VVPWL@0 tail gnd pwl (0ns 0 1.99ns 0 2ns 0.8 2.99ns 0.8 3ns 0) DC 0V AC 0V 0
VVPWL@1 head gnd pwl (0ps 0 0.99ns 0 1ns 0.8 1.99ns 0.8 2ns 0 2.99ns 0 3ns 0.8) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xcounter_@1 gnd head net_head0 net_head1 net_head2 net_head3 net_1 vdd net_16 tail net_tail0 net_tail1 net_tail2 net_tail3 net_0 ese370project2__counter_logic
.END
